** Profile: "SCHEMATIC1-sim6"  [ C:\EEC 111 Labs\Lab #6\Lab #6-PSpiceFiles\SCHEMATIC1\sim6.sim ] 

** Creating circuit file "sim6.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\EEC 111 Labs\Lab #6\Lab #6-PSpiceFiles\SCHEMATIC1\sim6\sim6_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\herob\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 2n 0 1p 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
