** Profile: "SCHEMATIC1-sim5"  [ C:\EEC 111 Labs\Lab #5\Lab #5-PSpiceFiles\SCHEMATIC1\sim5.sim ] 

** Creating circuit file "sim5.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\EEC 111 Labs\Lab #5\Lab #5-PSpiceFiles\SCHEMATIC1\sim5\sim5_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\herob\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_VIN 0 5 1m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
