** Profile: "SCHEMATIC1-sim4"  [ C:\EEC 111 Labs\Lab #4\Lab #4-PSpiceFiles\SCHEMATIC1\sim4.sim ] 

** Creating circuit file "sim4.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\EEC 111 Labs\Lab #4\Lab #4-PSpiceFiles\SCHEMATIC1\sim4\sim4_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\herob\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
